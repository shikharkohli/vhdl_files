library ieee;
use ieee.std_logic_1164.all;

entity mux2x1 is
    port(inp1,inp2:in std_logic;
         op(3 downto 0)
