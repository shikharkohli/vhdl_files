entity fulladder_tb is
end fulladder_tb;

architecture fulladder_tb_arch of fulladder_tb is
    component adder is
